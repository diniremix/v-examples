module main

fn main() {
	println('hola mundo en V')
	return
}
